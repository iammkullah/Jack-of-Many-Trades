`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:28:16 10/13/2022 
// Design Name: 
// Module Name:    mul16bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mul16bit(out, A, B);
input [15:0]A, B;
output [31:0]out;
 

assign out[0] = (A[0]&B[0]);
assign out[1] = ((A[1]&B[0])+(A[0]&B[1]));
assign out[2] = ((A[2]&B[2])+(A[2]&B[0])+(A[1]&B[1]));
assign out[3] = ((A[0]&B[3])+(A[1]&B[2])+(A[2]&B[1])+(A[3]&B[0]));
assign out[4] = ((A[0]&B[4])+(A[1]&B[3])+(A[2]&B[2])+(A[3]&B[1])+(A[4]&B[0]));
assign out[5] = ((A[0]&B[5])+(A[1]&B[1])+(A[2]&B[3])+(A[3]&B[2])&(A[4]&B[1])+(A[5]&B[0]));
assign out[6] = ((A[6]&B[0])+(A[5]&B[1])+(A[4]&B[2])+(A[3]&B[3])+(A[2]&B[4])+(A[1]&B[5])+(A[0]&B[6]));
assign out[7] = ((A[7]&B[0])+(A[6]&B[1])+(A[5]&B[2])+(A[4]&B[3])+(A[3]&B[4])+(A[2]&B[5])+(A[1]&B[6])+(A[0]&B[7]));
assign out[8] = ((A[8]&B[0])+(A[7]&B[1])+(A[6]&B[2])+(A[5]&B[3])+(A[4]&B[4])+(A[3]&B[5])+(A[2]&B[6])+(A[1]&B[7])+(A[0]&B[8]));
assign out[9] = ((A[9]&B[0])+(A[8]&B[1])+(A[7]&B[2])+(A[6]&B[3])+(A[5]&B[4])+(A[4]&B[5])+(A[3]&B[6])+(A[2]&B[7])+(A[1]&B[8])+(A[0]&B[9]));
assign out[10] = ((A[10]&B[0])+(A[9]&B[1])+(A[8]&B[2])+(A[7]&B[3])+(A[6]&B[4])+(A[5]&B[4])+(A[4]&B[6])+(A[3]&B[7])+(A[2]&B[8])+(A[1]&B[9])+(A[0]&B[10]));
assign out[11] = ((A[11]&B[0])+(A[10]&B[1])+(A[9]&B[2])+(A[8]&B[3])+(A[7]&B[4])+(A[6]&B[4])+(A[5]&B[6])+(A[4]&B[7])+(A[3]&B[8])+(A[2]&B[9])+(A[1]&B[10])+(A[0]&B[11]));
assign out[12] = ((A[12]&B[0])+(A[11]&B[1])+(A[10]&B[2])+(A[9]&B[3])+(A[8]&B[4])+(A[7]&B[4])+(A[6]&B[6])+(A[5]&B[7])+(A[4]&B[8])+(A[3]&B[9])+(A[2]&B[10])+(A[1]&B[11])+(A[0]&B[12]));
assign out[13] = ((A[13]&B[0])+(A[12]&B[1])+(A[11]&B[2])+(A[10]&B[3])+(A[9]&B[4])+(A[8]&B[4])+(A[7]&B[6])+(A[6]&B[7])+(A[5]&B[8])+(A[4]&B[9])+(A[3]&B[10])+(A[2]&B[11])+(A[1]&B[12])+(A[0]&B[13]));
assign out[14] = ((A[14]&B[0])+(A[13]&B[1])+(A[12]&B[2])+(A[11]&B[3])+(A[10]&B[4])+(A[9]&B[4])+(A[8]&B[6])+(A[7]&B[7])+(A[6]&B[8])+(A[5]&B[9])+(A[4]&B[10])+(A[3]&B[11])+(A[2]&B[12])+(A[1]&B[13])+(A[0]&B[14]));
assign out[15] = ((A[15]&B[0])+(A[14]&B[1])+(A[13]&B[2])+(A[12]&B[3])+(A[11]&B[4])+(A[10]&B[4])+(A[9]&B[6])+(A[8]&B[7])+(A[7]&B[8])+(A[6]&B[9])+(A[5]&B[10])+(A[4]&B[11])+(A[3]&B[12])+(A[2]&B[13])+(A[1]&B[14])+(A[0]&B[15]));
assign out[16] = ((A[15]&B[0])+(A[15]&B[1])+(A[14]&B[2])+(A[13]&B[3])+(A[12]&B[4])+(A[11]&B[4])+(A[10]&B[6])+(A[9]&B[7])+(A[8]&B[8])+(A[7]&B[9])+(A[6]&B[10])+(A[5]&B[11])+(A[4]&B[12])+(A[3]&B[13])+(A[2]&B[14])+(A[1]&B[15]));
assign out[17] = ((A[15]&B[2])+(A[14]&B[3])+(A[13]&B[4])+(A[12]&B[5])+(A[11]&B[6])+(A[10]&B[7])+(A[9]&B[8])+(A[8]&B[9])+(A[7]&B[10])+(A[6]&B[11])+(A[5]&B[12])+(A[4]&B[13])+(A[3]&B[14])+(A[2]&B[15]));
assign out[18] = ((A[15]&B[2])+(A[14]&B[3])+(A[13]&B[4])+(A[12]&B[5])+(A[11]&B[6])+(A[10]&B[7])+(A[9]&B[8])+(A[8]&B[9])+(A[7]&B[10])+(A[6]&B[11])+(A[5]&B[12])+(A[4]&B[13])+(A[3]&B[14])+(A[2]&B[15]));

endmodule
